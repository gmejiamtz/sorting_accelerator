
module ulx3s_sim (
    input clk_i,
    input reset_i,
    input a_i,
    input b_i,
    input c_i,
    output d_o 
);

top uut (.*);

endmodule
